`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:Ramya C
// Design Name: 1 bit Full adder
// Module Name: fa
//////////////////////////////////////////////////////////////////////////////////

module fa(a,b,cin,s,cout);
input a,b,cin;
output s,cout;
assign s=a^b^cin;
assign cout=(a&b)|(a&cin)|(b&cin);
endmodule
